-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
-- Created on Mon Sep 25 14:45:11 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY relogio IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        set : IN STD_LOGIC := '0';
        h_m : IN STD_LOGIC := '0';
        saida : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
    );
END relogio;

ARCHITECTURE BEHAVIOR OF relogio IS
    TYPE type_fstate IS (state1,horario,state2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,set,h_m)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= horario;
            saida <= "000";
        ELSE
            saida <= "000";
            CASE fstate IS
                WHEN state1 =>
                    IF (NOT((set = '1'))) THEN
                        reg_fstate <= horario;
                    ELSIF ((NOT((h_m = '1')) AND (set = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    saida <= "100";
                WHEN horario =>
                    IF (((set = '1') AND (h_m = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF (((set = '1') AND NOT((h_m = '1')))) THEN
                        reg_fstate <= state2;
                    ELSIF (NOT((set = '1'))) THEN
                        reg_fstate <= horario;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= horario;
                    END IF;

                    saida <= "001";
                WHEN state2 =>
                    IF (NOT((set = '1'))) THEN
                        reg_fstate <= horario;
                    ELSIF (((h_m = '1') AND (set = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    saida <= "010";
                WHEN OTHERS => 
                    saida <= "XXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
